module ADC_DCLK(CLR, RST_n,Enable, ADC_DCLK)

input CLR, RST_n,Enable;
output ADC_DCLK;


endmodule